module shift_right (
	IR,
	shift,
	B,
	H
);
	parameter data_length = 32;
	input IR;
	input [$clog2(data_length) - 1:0] shift;
	input [data_length - 1:0] B;
	output wire [data_length - 1:0] H;
	wire [($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)):($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length)] muxconnector;
	genvar i;
	genvar j;
	genvar k;
	generate
		for (j = 0; j < $clog2(data_length); j = j + 1) begin : genblk1
			for (i = 0; i < data_length; i = i + 1) begin : genblk1
				if ((i - (2 ** j)) >= 0) begin : genblk1
					mux_2to1 mx(
						.in_mux_x(muxconnector[(($clog2(data_length) >= 0 ? j : $clog2(data_length) - j) * data_length) + (i - (2 ** j))]),
						.in_mux_y(muxconnector[(($clog2(data_length) >= 0 ? j : $clog2(data_length) - j) * data_length) + i]),
						.s(shift[j]),
						.o_mux(muxconnector[(($clog2(data_length) >= 0 ? j + 1 : $clog2(data_length) - (j + 1)) * data_length) + i])
					);
				end
				else begin : genblk1
					mux_2to1 mx(
						.in_mux_x(IR),
						.in_mux_y(muxconnector[(($clog2(data_length) >= 0 ? j : $clog2(data_length) - j) * data_length) + i]),
						.s(shift[j]),
						.o_mux(muxconnector[(($clog2(data_length) >= 0 ? j + 1 : $clog2(data_length) - (j + 1)) * data_length) + i])
					);
				end
			end
		end
	endgenerate
	function automatic [(0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1:0] _sv2v_strm_10D6C;
		input reg [(0 + data_length) - 1:0] inp;
		reg [(0 + data_length) - 1:0] _sv2v_strm_55E18_inp;
		reg [(0 + data_length) - 1:0] _sv2v_strm_55E18_out;
		integer _sv2v_strm_55E18_idx;
		begin
			_sv2v_strm_55E18_inp = {inp};
			for (_sv2v_strm_55E18_idx = 0; _sv2v_strm_55E18_idx <= ((0 + data_length) - 1); _sv2v_strm_55E18_idx = _sv2v_strm_55E18_idx + 1)
				_sv2v_strm_55E18_out[((0 + data_length) - 1) - _sv2v_strm_55E18_idx-:1] = _sv2v_strm_55E18_inp[_sv2v_strm_55E18_idx+:1];
			_sv2v_strm_10D6C = ((0 + data_length) <= (0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) ? _sv2v_strm_55E18_out << ((0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - (0 + data_length)) : _sv2v_strm_55E18_out >> ((0 + data_length) - (0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length) + data_length) - 1)) + 1))));
		end
	endfunction
	assign {muxconnector[($clog2(data_length) >= 0 ? 0 : $clog2(data_length)) * data_length+:data_length]} = _sv2v_strm_10D6C({B});
	function automatic [data_length - 1:0] _sv2v_strm_AC36D;
		input reg [(0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1:0] inp;
		reg [(0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1:0] _sv2v_strm_55E18_inp;
		reg [(0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1:0] _sv2v_strm_55E18_out;
		integer _sv2v_strm_55E18_idx;
		begin
			_sv2v_strm_55E18_inp = {inp};
			for (_sv2v_strm_55E18_idx = 0; _sv2v_strm_55E18_idx <= ((0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1); _sv2v_strm_55E18_idx = _sv2v_strm_55E18_idx + 1)
				_sv2v_strm_55E18_out[((0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - 1) - _sv2v_strm_55E18_idx-:1] = _sv2v_strm_55E18_inp[_sv2v_strm_55E18_idx+:1];
			_sv2v_strm_AC36D = ((0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) <= data_length ? _sv2v_strm_55E18_out << (data_length - (0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1))) : _sv2v_strm_55E18_out >> ((0 + ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) >= (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) ? ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length)) + 1 : ((($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1 : ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) - (($clog2(data_length) >= 0 ? 0 : $clog2(data_length) * data_length) >= ($clog2(data_length) >= 0 ? (($clog2(data_length) + 1) * data_length) - 1 : ((1 - $clog2(data_length)) * data_length) + (($clog2(data_length) * data_length) - 1)) ? ($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length : ((($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length) + data_length) - 1)) + 1)) - data_length));
		end
	endfunction
	assign H = _sv2v_strm_AC36D({muxconnector[($clog2(data_length) >= 0 ? $clog2(data_length) : $clog2(data_length) - $clog2(data_length)) * data_length+:data_length]});
endmodule
